//********************************************************************                                        
//  AUTHOR: Engineering Design Institute/ASIC Design and Verification	                                                     		
//  DESCRIPTION: Arbiter Interface                                        
//  MODULE NAME: arb_if
//********************************************************************
 `timescale 10 ns / 1 ps

 interface arb_if(input bit clk);
	logic [1:0] grant, request;
	logic reset;
 endinterface

 

 
 
 

 
 
 
 
 