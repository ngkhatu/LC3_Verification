class Assertions

endclass

