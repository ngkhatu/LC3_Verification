
class Monitor

endclass
