
class Agent

endclass

