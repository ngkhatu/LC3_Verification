class Checker

endclass
