library verilog;
use verilog.vl_types.all;
entity dut_Probe_if is
    port(
        fetch_enable_updatePC: in     vl_logic;
        fetch_enable_fetch: in     vl_logic;
        fetch_br_taken  : in     vl_logic;
        fetch_taddr     : in     vl_logic_vector(15 downto 0);
        fetch_instrmem_rd: in     vl_logic;
        fetch_pc        : in     vl_logic_vector(15 downto 0);
        fetch_npc_out   : in     vl_logic_vector(15 downto 0);
        decode_enable_decode: in     vl_logic;
        decode_Instr_dout: in     vl_logic_vector(15 downto 0);
        decode_npc_out  : in     vl_logic_vector(15 downto 0);
        decode_IR       : in     vl_logic_vector(15 downto 0);
        decode_npc_in   : in     vl_logic_vector(15 downto 0);
        decode_Mem_control: in     vl_logic;
        decode_E_control: in     vl_logic_vector(5 downto 0);
        decode_W_control: in     vl_logic_vector(1 downto 0);
        control_IR      : in     vl_logic_vector(15 downto 0);
        control_IR_Exec : in     vl_logic_vector(15 downto 0);
        control_IMem_dout: in     vl_logic_vector(15 downto 0);
        control_complete_data: in     vl_logic;
        control_complete_instr: in     vl_logic;
        control_nzp     : in     vl_logic_vector(2 downto 0);
        control_psr     : in     vl_logic_vector(2 downto 0);
        control_enable_fetch: in     vl_logic;
        control_enable_updatePC: in     vl_logic;
        control_enable_decode: in     vl_logic;
        control_enable_execute: in     vl_logic;
        control_enable_writeback: in     vl_logic;
        control_br_taken: in     vl_logic;
        control_bypass_alu_1: in     vl_logic;
        control_bypass_alu_2: in     vl_logic;
        control_bypass_mem_1: in     vl_logic;
        control_bypass_mem_2: in     vl_logic;
        control_mem_state: in     vl_logic_vector(1 downto 0);
        ex_E_control    : in     vl_logic_vector(5 downto 0);
        ex_IR           : in     vl_logic_vector(15 downto 0);
        ex_npc_in       : in     vl_logic_vector(15 downto 0);
        ex_VSR1         : in     vl_logic_vector(15 downto 0);
        ex_VSR2         : in     vl_logic_vector(15 downto 0);
        ex_bypass_alu_1 : in     vl_logic;
        ex_bypass_alu_2 : in     vl_logic;
        ex_bypass_mem_1 : in     vl_logic;
        ex_bypass_mem_2 : in     vl_logic;
        ex_Mem_control_in: in     vl_logic;
        ex_Mem_control_out: in     vl_logic;
        ex_enable_execute: in     vl_logic;
        ex_W_Control_in : in     vl_logic_vector(1 downto 0);
        ex_W_Control_out: in     vl_logic_vector(1 downto 0);
        ex_Mem_bypass_value: in     vl_logic_vector(15 downto 0);
        ex_M_data       : in     vl_logic_vector(15 downto 0);
        ex_IR_exec      : in     vl_logic_vector(15 downto 0);
        ex_aluout       : in     vl_logic_vector(15 downto 0);
        ex_pcout        : in     vl_logic_vector(15 downto 0);
        ex_dr           : in     vl_logic_vector(2 downto 0);
        ex_sr1          : in     vl_logic_vector(2 downto 0);
        ex_sr2          : in     vl_logic_vector(2 downto 0);
        ex_NZP          : in     vl_logic_vector(2 downto 0);
        execute_pcout   : in     vl_logic_vector(15 downto 0);
        writeback_enable_writeback: in     vl_logic;
        writeback_sr1   : in     vl_logic_vector(2 downto 0);
        writeback_sr2   : in     vl_logic_vector(2 downto 0);
        writeback_dr    : in     vl_logic_vector(2 downto 0);
        writeback_psr   : in     vl_logic_vector(2 downto 0);
        writeback_aluout: in     vl_logic_vector(15 downto 0);
        writeback_memout: in     vl_logic_vector(15 downto 0);
        writeback_pcout : in     vl_logic_vector(15 downto 0);
        writeback_VSR1  : in     vl_logic_vector(15 downto 0);
        writeback_VSR2  : in     vl_logic_vector(15 downto 0);
        wr_R0           : in     vl_logic_vector(15 downto 0);
        wr_R1           : in     vl_logic_vector(15 downto 0);
        wr_R2           : in     vl_logic_vector(15 downto 0);
        wr_R3           : in     vl_logic_vector(15 downto 0);
        wr_R4           : in     vl_logic_vector(15 downto 0);
        wr_R5           : in     vl_logic_vector(15 downto 0);
        wr_R6           : in     vl_logic_vector(15 downto 0);
        wr_R7           : in     vl_logic_vector(15 downto 0);
        MemAccess_M_Data: in     vl_logic_vector(15 downto 0);
        MemAccess_M_Addr: in     vl_logic_vector(15 downto 0);
        MemAccess_DMem_dout: in     vl_logic_vector(15 downto 0);
        MemAccess_DMem_addr: in     vl_logic_vector(15 downto 0);
        MemAccess_DMem_din: in     vl_logic_vector(15 downto 0);
        MemAccess_DMem_rd: in     vl_logic;
        MemAccess_M_Control: in     vl_logic;
        MemAccess_mem_state: in     vl_logic_vector(1 downto 0);
        writeback_W_control: in     vl_logic_vector(1 downto 0)
    );
end dut_Probe_if;
