library verilog;
use verilog.vl_types.all;
entity data_def_test_v_unit is
end data_def_test_v_unit;
