library verilog;
use verilog.vl_types.all;
entity Instruction_sv_unit is
end Instruction_sv_unit;
