library verilog;
use verilog.vl_types.all;
entity LC3_test_top is
    generic(
        simulation_cycle: integer := 20
    );
end LC3_test_top;
